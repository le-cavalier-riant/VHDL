library ieee;
use ieee.std_logic_1164.all;

entity module is
	port (horloge: in std_logic);
end module;

architecture Behavioral of module is begin end Behavioral;